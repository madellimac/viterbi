
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package definition_pkg is
 
    type state_metric_array is array(0 to 7) of std_logic_vector(6 downto 0);
	 type branch_metric_array is array(0 to 3) of std_logic_vector(3 downto 0);

end definition_pkg;

package body definition_pkg is

 
end definition_pkg;
